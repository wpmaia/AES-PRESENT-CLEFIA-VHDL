----------------------------------------------------------------------------------
-- Mestrado em Engenharia El�trica (Universidade Federal de Sergipe UFS - Brasil)
-- Disserta��o: Projeto, Implementa��o e Desempenho dos Algoritmos Criptogr�ficos
-- AES, PRESENT e CLEFIA em FPGA
-- Autor: William Pedrosa Maia
-- E-mail: wmaia.eng@gmail.com
-- Prof. Orientador: Edward David Moreno
-- Data: Julho/2017
--
-- Projeto: CLEFIA-128                                                                                                                                                                                       
--
-- Descri��o: S1 (Tabela de Substitui��o S1)
-- Vers�o: 1
--                                                                                                                                                      
-- Adaptado de (Sony Corporation, 2010)                                                                                    
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity S1 is
    Port ( s1_in : in STD_LOGIC_VECTOR (7 downto 0);
           s1_out : out STD_LOGIC_VECTOR (7 downto 0)
           );
end S1;

architecture Behavioral of S1 is

begin

	 with s1_in  (7 downto 0) select
          s1_out (7 downto 0) <=
         
		  "01101100"	when	"00000000",	--(X"6c")	0
          "11011010"	when	"00000001",	--(X"da")	1
          "11000011"	when	"00000010",	--(X"c3")	2
          "11101001"	when	"00000011",	--(X"e9")	3
          "01001110"	when	"00000100",	--(X"4e")	4
          "10011101"	when	"00000101",	--(X"9d")	5
          "00001010"	when	"00000110",	--(X"0a")	6
          "00111101"	when	"00000111",	--(X"3d")	7
          "10111000"	when	"00001000",	--(X"b8")	8
          "00110110"	when	"00001001",	--(X"36")	9
          "10110100"	when	"00001010",	--(X"b4")	10
          "00111000"	when	"00001011",	--(X"38")	11
          "00010011"	when	"00001100",	--(X"13")	12
          "00110100"	when	"00001101",	--(X"34")	13
          "00001100"	when	"00001110",	--(X"0c")	14
          "11011001"	when	"00001111",	--(X"d9")	15
          "10111111"	when	"00010000",	--(X"bf")	16
          "01110100"	when	"00010001",	--(X"74")	17
          "10010100"	when	"00010010",	--(X"94")	18
          "10001111"	when	"00010011",	--(X"8f")	19
          "10110111"	when	"00010100",	--(X"b7")	20
          "10011100"	when	"00010101",	--(X"9c")	21
          "11100101"	when	"00010110",	--(X"e5")	22
          "11011100"	when	"00010111",	--(X"dc")	23
          "10011110"	when	"00011000",	--(X"9e")	24
          "00000111"	when	"00011001",	--(X"7")	25
          "01001001"	when	"00011010",	--(X"49")	26
          "01001111"	when	"00011011",	--(X"4f")	27
          "10011000"	when	"00011100",	--(X"98")	28
          "00101100"	when	"00011101",	--(X"2c")	29
          "10110000"	when	"00011110",	--(X"b0")	30
          "10010011"	when	"00011111",	--(X"93")	31
          "00010010"	when	"00100000",	--(X"12")	32
          "11101011"	when	"00100001",	--(X"eb")	33
          "11001101"	when	"00100010",	--(X"cd")	34
          "10110011"	when	"00100011",	--(X"b3")	35
          "10010010"	when	"00100100",	--(X"92")	36
          "11100111"	when	"00100101",	--(X"e7")	37
          "01000001"	when	"00100110",	--(X"41")	38
          "01100000"	when	"00100111",	--(X"60")	39
          "11100011"	when	"00101000",	--(X"e3")	40
          "00100001"	when	"00101001",	--(X"21")	41
          "00100111"	when	"00101010",	--(X"27")	42
          "00111011"	when	"00101011",	--(X"3b")	43
          "11100110"	when	"00101100",	--(X"e6")	44
          "00011001"	when	"00101101",	--(X"19")	45
          "11010010"	when	"00101110",	--(X"d2")	46
          "00001110"	when	"00101111",	--(X"0e")	47
          "10010001"	when	"00110000",	--(X"91")	48
          "00010001"	when	"00110001",	--(X"11")	49
          "11000111"	when	"00110010",	--(X"c7")	50
          "00111111"	when	"00110011",	--(X"3f")	51
          "00101010"	when	"00110100",	--(X"2a")	52
          "10001110"	when	"00110101",	--(X"8e")	53
          "10100001"	when	"00110110",	--(X"a1")	54
          "10111100"	when	"00110111",	--(X"bc")	55
          "00101011"	when	"00111000",	--(X"2b")	56
          "11001000"	when	"00111001",	--(X"c8")	57
          "11000101"	when	"00111010",	--(X"c5")	58
          "00001111"	when	"00111011",	--(X"0f")	59
          "01011011"	when	"00111100",	--(X"5b")	60
          "11110011"	when	"00111101",	--(X"f3")	61
          "10000111"	when	"00111110",	--(X"87")	62
          "10001011"	when	"00111111",	--(X"8b")	63
          "11111011"	when	"01000000",	--(X"fb")	64
          "11110101"	when	"01000001",	--(X"f5")	65
          "11011110"	when	"01000010",	--(X"de")	66
          "00100000"	when	"01000011",	--(X"20")	67
          "11000110"	when	"01000100",	--(X"c6")	68
          "10100111"	when	"01000101",	--(X"a7")	69
          "10000100"	when	"01000110",	--(X"84")	70
          "11001110"	when	"01000111",	--(X"ce")	71
          "11011000"	when	"01001000",	--(X"d8")	72
          "01100101"	when	"01001001",	--(X"65")	73
          "01010001"	when	"01001010",	--(X"51")	74
          "11001001"	when	"01001011",	--(X"c9")	75
          "10100100"	when	"01001100",	--(X"a4")	76
          "11101111"	when	"01001101",	--(X"ef")	77
          "01000011"	when	"01001110",	--(X"43")	78
          "01010011"	when	"01001111",	--(X"53")	79
          "00100101"	when	"01010000",	--(X"25")	80
          "01011101"	when	"01010001",	--(X"5d")	81
          "10011011"	when	"01010010",	--(X"9b")	82
          "00110001"	when	"01010011",	--(X"31")	83
          "11101000"	when	"01010100",	--(X"e8")	84
          "00111110"	when	"01010101",	--(X"3e")	85
          "00001101"	when	"01010110",	--(X"0d")	86
          "11010111"	when	"01010111",	--(X"d7")	87
          "10000000"	when	"01011000",	--(X"80")	88
          "11111111"	when	"01011001",	--(X"ff")	89
          "01101001"	when	"01011010",	--(X"69")	90
          "10001010"	when	"01011011",	--(X"8a")	91
          "10111010"	when	"01011100",	--(X"ba")	92
          "00001011"	when	"01011101",	--(X"0b")	93
          "01110011"	when	"01011110",	--(X"73")	94
          "01011100"	when	"01011111",	--(X"5c")	95
          "01101110"	when	"01100000",	--(X"6e")	96
          "01010100"	when	"01100001",	--(X"54")	97
          "00010101"	when	"01100010",	--(X"15")	98
          "01100010"	when	"01100011",	--(X"62")	99
          "11110110"	when	"01100100",	--(X"f6")	100
          "00110101"	when	"01100101",	--(X"35")	101
          "00110000"	when	"01100110",	--(X"30")	102
          "01010010"	when	"01100111",	--(X"52")	103
          "10100011"	when	"01101000",	--(X"a3")	104
          "00010110"	when	"01101001",	--(X"16")	105
          "11010011"	when	"01101010",	--(X"d3")	106
          "00101000"	when	"01101011",	--(X"28")	107
          "00110010"	when	"01101100",	--(X"32")	108
          "11111010"	when	"01101101",	--(X"fa")	109
          "10101010"	when	"01101110",	--(X"aa")	110
          "01011110"	when	"01101111",	--(X"5e")	111
          "11001111"	when	"01110000",	--(X"cf")	112
          "11101010"	when	"01110001",	--(X"ea")	113
          "11101101"	when	"01110010",	--(X"ed")	114
          "01111000"	when	"01110011",	--(X"78")	115
          "00110011"	when	"01110100",	--(X"33")	116
          "01011000"	when	"01110101",	--(X"58")	117
          "00001001"	when	"01110110",	--(X"9")	118
          "01111011"	when	"01110111",	--(X"7b")	119
          "01100011"	when	"01111000",	--(X"63")	120
          "11000000"	when	"01111001",	--(X"c0")	121
          "11000001"	when	"01111010",	--(X"c1")	122
          "01000110"	when	"01111011",	--(X"46")	123
          "00011110"	when	"01111100",	--(X"1e")	124
          "11011111"	when	"01111101",	--(X"df")	125
          "10101001"	when	"01111110",	--(X"a9")	126
          "10011001"	when	"01111111",	--(X"99")	127
          "01010101"	when	"10000000",	--(X"55")	128
          "00000100"	when	"10000001",	--(X"4")	129
          "11000100"	when	"10000010",	--(X"c4")	130
          "10000110"	when	"10000011",	--(X"86")	131
          "00111001"	when	"10000100",	--(X"39")	132
          "01110111"	when	"10000101",	--(X"77")	133
          "10000010"	when	"10000110",	--(X"82")	134
          "11101100"	when	"10000111",	--(X"ec")	135
          "01000000"	when	"10001000",	--(X"40")	136
          "00011000"	when	"10001001",	--(X"18")	137
          "10010000"	when	"10001010",	--(X"90")	138
          "10010111"	when	"10001011",	--(X"97")	139
          "01011001"	when	"10001100",	--(X"59")	140
          "11011101"	when	"10001101",	--(X"dd")	141
          "10000011"	when	"10001110",	--(X"83")	142
          "00011111"	when	"10001111",	--(X"1f")	143
          "10011010"	when	"10010000",	--(X"9a")	144
          "00110111"	when	"10010001",	--(X"37")	145
          "00000110"	when	"10010010",	--(X"6")	146
          "00100100"	when	"10010011",	--(X"24")	147
          "01100100"	when	"10010100",	--(X"64")	148
          "01111100"	when	"10010101",	--(X"7c")	149
          "10100101"	when	"10010110",	--(X"a5")	150
          "01010110"	when	"10010111",	--(X"56")	151
          "01001000"	when	"10011000",	--(X"48")	152
          "00001000"	when	"10011001",	--(X"8")	153
          "10000101"	when	"10011010",	--(X"85")	154
          "11010000"	when	"10011011",	--(X"d0")	155
          "01100001"	when	"10011100",	--(X"61")	156
          "00100110"	when	"10011101",	--(X"26")	157
          "11001010"	when	"10011110",	--(X"ca")	158
          "01101111"	when	"10011111",	--(X"6f")	159
          "01111110"	when	"10100000",	--(X"7e")	160
          "01101010"	when	"10100001",	--(X"6a")	161
          "10110110"	when	"10100010",	--(X"b6")	162
          "01110001"	when	"10100011",	--(X"71")	163
          "10100000"	when	"10100100",	--(X"a0")	164
          "01110000"	when	"10100101",	--(X"70")	165
          "00000101"	when	"10100110",	--(X"5")	166
          "11010001"	when	"10100111",	--(X"d1")	167
          "01000101"	when	"10101000",	--(X"45")	168
          "10001100"	when	"10101001",	--(X"8c")	169
          "00100011"	when	"10101010",	--(X"23")	170
          "00011100"	when	"10101011",	--(X"1c")	171
          "11110000"	when	"10101100",	--(X"f0")	172
          "11101110"	when	"10101101",	--(X"ee")	173
          "10001001"	when	"10101110",	--(X"89")	174
          "10101101"	when	"10101111",	--(X"ad")	175
          "01111010"	when	"10110000",	--(X"7a")	176
          "01001011"	when	"10110001",	--(X"4b")	177
          "11000010"	when	"10110010",	--(X"c2")	178
          "00101111"	when	"10110011",	--(X"2f")	179
          "11011011"	when	"10110100",	--(X"db")	180
          "01011010"	when	"10110101",	--(X"5a")	181
          "01001101"	when	"10110110",	--(X"4d")	182
          "01110110"	when	"10110111",	--(X"76")	183
          "01100111"	when	"10111000",	--(X"67")	184
          "00010111"	when	"10111001",	--(X"17")	185
          "00101101"	when	"10111010",	--(X"2d")	186
          "11110100"	when	"10111011",	--(X"f4")	187
          "11001011"	when	"10111100",	--(X"cb")	188
          "10110001"	when	"10111101",	--(X"b1")	189
          "01001010"	when	"10111110",	--(X"4a")	190
          "10101000"	when	"10111111",	--(X"a8")	191
          "10110101"	when	"11000000",	--(X"b5")	192
          "00100010"	when	"11000001",	--(X"22")	193
          "01000111"	when	"11000010",	--(X"47")	194
          "00111010"	when	"11000011",	--(X"3a")	195
          "11010101"	when	"11000100",	--(X"d5")	196
          "00010000"	when	"11000101",	--(X"10")	197
          "01001100"	when	"11000110",	--(X"4c")	198
          "01110010"	when	"11000111",	--(X"72")	199
          "11001100"	when	"11001000",	--(X"cc")	200
          "00000000"	when	"11001001",	--(X"0")	201
          "11111001"	when	"11001010",	--(X"f9")	202
          "11100000"	when	"11001011",	--(X"e0")	203
          "11111101"	when	"11001100",	--(X"fd")	204
          "11100010"	when	"11001101",	--(X"e2")	205
          "11111110"	when	"11001110",	--(X"fe")	206
          "10101110"	when	"11001111",	--(X"ae")	207
          "11111000"	when	"11010000",	--(X"f8")	208
          "01011111"	when	"11010001",	--(X"5f")	209
          "10101011"	when	"11010010",	--(X"ab")	210
          "11110001"	when	"11010011",	--(X"f1")	211
          "00011011"	when	"11010100",	--(X"1b")	212
          "01000010"	when	"11010101",	--(X"42")	213
          "10000001"	when	"11010110",	--(X"81")	214
          "11010110"	when	"11010111",	--(X"d6")	215
          "10111110"	when	"11011000",	--(X"be")	216
          "01000100"	when	"11011001",	--(X"44")	217
          "00101001"	when	"11011010",	--(X"29")	218
          "10100110"	when	"11011011",	--(X"a6")	219
          "01010111"	when	"11011100",	--(X"57")	220
          "10111001"	when	"11011101",	--(X"b9")	221
          "10101111"	when	"11011110",	--(X"af")	222
          "11110010"	when	"11011111",	--(X"f2")	223
          "11010100"	when	"11100000",	--(X"d4")	224
          "01110101"	when	"11100001",	--(X"75")	225
          "01100110"	when	"11100010",	--(X"66")	226
          "10111011"	when	"11100011",	--(X"bb")	227
          "01101000"	when	"11100100",	--(X"68")	228
          "10011111"	when	"11100101",	--(X"9f")	229
          "01010000"	when	"11100110",	--(X"50")	230
          "00000010"	when	"11100111",	--(X"2")	231
          "00000001"	when	"11101000",	--(X"1")	232
          "00111100"	when	"11101001",	--(X"3c")	233
          "01111111"	when	"11101010",	--(X"7f")	234
          "10001101"	when	"11101011",	--(X"8d")	235
          "00011010"	when	"11101100",	--(X"1a")	236
          "10001000"	when	"11101101",	--(X"88")	237
          "10111101"	when	"11101110",	--(X"bd")	238
          "10101100"	when	"11101111",	--(X"ac")	239
          "11110111"	when	"11110000",	--(X"f7")	240
          "11100100"	when	"11110001",	--(X"e4")	241
          "01111001"	when	"11110010",	--(X"79")	242
          "10010110"	when	"11110011",	--(X"96")	243
          "10100010"	when	"11110100",	--(X"a2")	244
          "11111100"	when	"11110101",	--(X"fc")	245
          "01101101"	when	"11110110",	--(X"6d")	246
          "10110010"	when	"11110111",	--(X"b2")	247
          "01101011"	when	"11111000",	--(X"6b")	248
          "00000011"	when	"11111001",	--(X"3")	249
          "11100001"	when	"11111010",	--(X"e1")	250
          "00101110"	when	"11111011",	--(X"2e")	251
          "01111101"	when	"11111100",	--(X"7d")	252
          "00010100"	when	"11111101",	--(X"14")	253
          "10010101"	when	"11111110",	--(X"95")	254
          "00011101"	when	"11111111",	--(X"1d")	255        
                                                         
         "XXXXXXXX" WHEN OTHERS;

end Behavioral;
