----------------------------------------------------------------------------------
-- Mestrado em Engenharia El�trica (Universidade Federal de Sergipe UFS - Brasil)
-- Disserta��o: Projeto, Implementa��o e Desempenho dos Algoritmos Criptogr�ficos
-- AES, PRESENT e CLEFIA em FPGA
-- Autor: William Pedrosa Maia
-- E-mail: wmaia.eng@gmail.com
-- Prof. Orientador: Edward David Moreno
-- Data: Julho/2017
--
-- Projeto: CLEFIA-128                                                                                                                                                                                       
--
-- Descri��o: Constants (Constantes predefinidas para a gera��o das subchaves)
-- Vers�o: 1
--                                                                                                                                                      
-- Adaptado de (Sony Corporation, 2010)                                                                                    
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity const is
 	Port (
 	 	  clk     : in std_logic;
 	 	  reset   : in std_logic;
 	 	  enable  : in std_logic;
 	 	  const_l : out std_logic_vector (63 downto 0)
 	 	  );
end const;

architecture Behavioral of const is
	
	signal sig_const : std_logic_vector (63 downto 0) := (others => '0');
	type memory is array (1 to 60) of std_logic_vector(31 downto 0);
	constant myrom : memory := (
-- Constants Key Shedule (for 128-bit key)
1 => "11110101011010110111101011101011", --f56b7aeb
2  => "10011001010010101000101001000010", --994a8a42
3  => "10010110101001001011110101110101", --96a4bd75
4  => "11111010100001010100010100100001", --fa854521
5  => "01110011010110110111011010001010", --735b768a
6  => "00011111011110101011101011000100", --1f7abac4
7  => "11010101101111000011101101000101", --d5bc3b45
8  => "10111001100111010101110101100010", --b99d5d62
9  => "01010010110101110011010110010010", --52d73592
10 => "00111110111101100011011011100101", --3ef636e5
11 => "11000101011110100001101011001001", --c57a1ac9
12 => "10101001010110111001101101110010", --a95b9b72
13 => "01011010101101000010010101010100", --5ab42554
14 => "00110110100101010101010111101101", --369555ed
15 => "00010101010100111011101010011010", --1553ba9a
16 => "01111001011100101011001010100010", --7972b2a2
17 => "11100110101110000101110101001101", --e6b85d4d
18 => "10001010100110010101100101010001", --8a995951
19 => "01001011010101010000011010010110", --4b550696
20 => "00100111011101001011010011111100", --2774b4fc
21 => "11001001101110110000001101001011", --c9bb034b
22 => "10100101100110100101101001111110", --a59a5a7e
23 => "10001000110011001000000110100101", --88cc81a5
24 => "11100100111011010010110100111111", --e4ed2d3f
25 => "01111100011011110110100011100010", --7c6f68e2
26 => "00010000010011101000111011001011", --104e8ecb
27 => "11010010001001100011010001110001", --d2263471
28 => "10111110000001111100011101100101", --be07c765
29 => "01010001000110100011001000001000", --511a3208
30 => "00111101001110111111101111100110", --3d3bfbe6
31 => "00010000100001001011000100110100", --1084b134
32 => "01111100101001010110010110100111", --7ca565a7
33 => "00110000010010111111000010101010", --304bf0aa
34 => "01011100011010101010101010000111", --5c6aaa87
35 => "11110100001101000111100001010101", --f4347855
36 => "10011000000101011101010101000011", --9815d543
37 => "01000010000100110001010000011010", --4213141a
38 => "00101110001100101111001011110101", --2e32f2f5
39 => "11001101000110000000101000001101", --cd180a0d
40 => "10100001001110011111100101111010", --a139f97a
41 => "01011110100001010010110100110110", --5e852d36
42 => "00110010101001000110010011101001", --32a464e9
43 => "11000011010100110001011010011011", --c353169b
44 => "10101111011100101011001001110100", --af72b274
45 => "10001101101110001000101101001101", --8db88b4d
46 => "11100001100110010101100100111010", --e199593a
47 => "01111110110101010110110110010110", --7ed56d96
48 => "00010010111101000011010011001001", --12f434c9
49 => "11010011011110110011011011001011", --d37b36cb
50 => "10111111010110101001101001100100", --bf5a9a64
51 => "10000101101011001001101101100101", --85ac9b65
52 => "11101001100011010100110100110010", --e98d4d32
53 => "01111010110111110110010110000010", --7adf6582
54 => "00010110111111100011111011001101", --16fe3ecd
55 => "11010001011111100011001011000001", --d17e32c1
56 => "10111101010111111001111101100110", --bd5f9f66
57 => "01010000101101100011000101010000", --50b63150
58 => "00111100100101110101011111100111", --3c9757e7
59 => "00010000010100101011000010011000", --1052b098
60 => "01111100011100111011001110100111", --7c73b3a7
others => "00000000000000000000000000000000");

begin
	
	key_const : process (clk, reset, enable)
	variable internal_count : integer range 0 to 30;	
		begin
			if (reset = '1') then
				internal_count := 0;
				sig_const  <= (others => '0');
			elsif (clk = '1' and clk'Event) then
				if (enable = '1') then	 
				internal_count := internal_count + 1;
				sig_const <= myrom((internal_count*2)-1) & myrom(internal_count*2);
				if (internal_count = 30) then                        
				    internal_count := 0;
					end if;
				end if;
			end if;
		end process key_const;	
	
const_l  <= sig_const;

end Behavioral;