----------------------------------------------------------------------------------
-- Mestrado em Engenharia El�trica (Universidade Federal de Sergipe UFS - Brasil)
-- Disserta��o: Projeto, Implementa��o e Desempenho dos Algoritmos Criptogr�ficos
-- AES, PRESENT e CLEFIA em FPGA
-- Autor: William Pedrosa Maia
-- E-mail: wmaia.eng@gmail.com
-- Prof. Orientador: Edward David Moreno
-- Data: Julho/2017
--
-- Projeto: CLEFIA-128                                                                                                                                                                                       
--
-- Descri��o: S0 (Tabela de Substitui��o S0)
-- Vers�o: 1
--                                                                                                                                                      
-- Adaptado de (Sony Corporation, 2010)                                                                                    
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity S0 is
    Port ( s0_in : in STD_LOGIC_VECTOR (7 downto 0);
           s0_out : out STD_LOGIC_VECTOR (7 downto 0)
           );
end S0;

architecture Behavioral of S0 is

begin

	 with s0_in  (7 downto 0) select
          s0_out (7 downto 0) <=
         
		  "01010111"	when	"00000000",	--(X"57")	0
          "01001001"	when	"00000001",	--(X"49")	1
          "11010001"	when	"00000010",	--(X"d1")	2
          "11000110"	when	"00000011",	--(X"c6")	3
          "00101111"	when	"00000100",	--(X"2f")	4
          "00110011"	when	"00000101",	--(X"33")	5
          "01110100"	when	"00000110",	--(X"74")	6
          "11111011"	when	"00000111",	--(X"fb")	7
          "10010101"	when	"00001000",	--(X"95")	8
          "01101101"	when	"00001001",	--(X"6d")	9
          "10000010"	when	"00001010",	--(X"82")	10
          "11101010"	when	"00001011",	--(X"ea")	11
          "00001110"	when	"00001100",	--(X"0e")	12
          "10110000"	when	"00001101",	--(X"b0")	13
          "10101000"	when	"00001110",	--(X"a8")	14
          "00011100"	when	"00001111",	--(X"1c")	15
          "00101000"	when	"00010000",	--(X"28")	16
          "11010000"	when	"00010001",	--(X"d0")	17
          "01001011"	when	"00010010",	--(X"4b")	18
          "10010010"	when	"00010011",	--(X"92")	19
          "01011100"	when	"00010100",	--(X"5c")	20
          "11101110"	when	"00010101",	--(X"ee")	21
          "10000101"	when	"00010110",	--(X"85")	22
          "10110001"	when	"00010111",	--(X"b1")	23
          "11000100"	when	"00011000",	--(X"c4")	24
          "00001010"	when	"00011001",	--(X"0a")	25
          "01110110"	when	"00011010",	--(X"76")	26
          "00111101"	when	"00011011",	--(X"3d")	27
          "01100011"	when	"00011100",	--(X"63")	28
          "11111001"	when	"00011101",	--(X"f9")	29
          "00010111"	when	"00011110",	--(X"17")	30
          "10101111"	when	"00011111",	--(X"af")	31
          "10111111"	when	"00100000",	--(X"bf")	32
          "10100001"	when	"00100001",	--(X"a1")	33
          "00011001"	when	"00100010",	--(X"19")	34
          "01100101"	when	"00100011",	--(X"65")	35
          "11110111"	when	"00100100",	--(X"f7")	36
          "01111010"	when	"00100101",	--(X"7a")	37
          "00110010"	when	"00100110",	--(X"32")	38
          "00100000"	when	"00100111",	--(X"20")	39
          "00000110"	when	"00101000",	--(X"6")	40
          "11001110"	when	"00101001",	--(X"ce")	41
          "11100100"	when	"00101010",	--(X"e4")	42
          "10000011"	when	"00101011",	--(X"83")	43
          "10011101"	when	"00101100",	--(X"9d")	44
          "01011011"	when	"00101101",	--(X"5b")	45
          "01001100"	when	"00101110",	--(X"4c")	46
          "11011000"	when	"00101111",	--(X"d8")	47
          "01000010"	when	"00110000",	--(X"42")	48
          "01011101"	when	"00110001",	--(X"5d")	49
          "00101110"	when	"00110010",	--(X"2e")	50
          "11101000"	when	"00110011",	--(X"e8")	51
          "11010100"	when	"00110100",	--(X"d4")	52
          "10011011"	when	"00110101",	--(X"9b")	53
          "00001111"	when	"00110110",	--(X"0f")	54
          "00010011"	when	"00110111",	--(X"13")	55
          "00111100"	when	"00111000",	--(X"3c")	56
          "10001001"	when	"00111001",	--(X"89")	57
          "01100111"	when	"00111010",	--(X"67")	58
          "11000000"	when	"00111011",	--(X"c0")	59
          "01110001"	when	"00111100",	--(X"71")	60
          "10101010"	when	"00111101",	--(X"aa")	61
          "10110110"	when	"00111110",	--(X"b6")	62
          "11110101"	when	"00111111",	--(X"f5")	63
          "10100100"	when	"01000000",	--(X"a4")	64
          "10111110"	when	"01000001",	--(X"be")	65
          "11111101"	when	"01000010",	--(X"fd")	66
          "10001100"	when	"01000011",	--(X"8c")	67
          "00010010"	when	"01000100",	--(X"12")	68
          "00000000"	when	"01000101",	--(X"0")	69
          "10010111"	when	"01000110",	--(X"97")	70
          "11011010"	when	"01000111",	--(X"da")	71
          "01111000"	when	"01001000",	--(X"78")	72
          "11100001"	when	"01001001",	--(X"e1")	73
          "11001111"	when	"01001010",	--(X"cf")	74
          "01101011"	when	"01001011",	--(X"6b")	75
          "00111001"	when	"01001100",	--(X"39")	76
          "01000011"	when	"01001101",	--(X"43")	77
          "01010101"	when	"01001110",	--(X"55")	78
          "00100110"	when	"01001111",	--(X"26")	79
          "00110000"	when	"01010000",	--(X"30")	80
          "10011000"	when	"01010001",	--(X"98")	81
          "11001100"	when	"01010010",	--(X"cc")	82
          "11011101"	when	"01010011",	--(X"dd")	83
          "11101011"	when	"01010100",	--(X"eb")	84
          "01010100"	when	"01010101",	--(X"54")	85
          "10110011"	when	"01010110",	--(X"b3")	86
          "10001111"	when	"01010111",	--(X"8f")	87
          "01001110"	when	"01011000",	--(X"4e")	88
          "00010110"	when	"01011001",	--(X"16")	89
          "11111010"	when	"01011010",	--(X"fa")	90
          "00100010"	when	"01011011",	--(X"22")	91
          "10100101"	when	"01011100",	--(X"a5")	92
          "01110111"	when	"01011101",	--(X"77")	93
          "00001001"	when	"01011110",	--(X"9")	94
          "01100001"	when	"01011111",	--(X"61")	95
          "11010110"	when	"01100000",	--(X"d6")	96
          "00101010"	when	"01100001",	--(X"2a")	97
          "01010011"	when	"01100010",	--(X"53")	98
          "00110111"	when	"01100011",	--(X"37")	99
          "01000101"	when	"01100100",	--(X"45")	100
          "11000001"	when	"01100101",	--(X"c1")	101
          "01101100"	when	"01100110",	--(X"6c")	102
          "10101110"	when	"01100111",	--(X"ae")	103
          "11101111"	when	"01101000",	--(X"ef")	104
          "01110000"	when	"01101001",	--(X"70")	105
          "00001000"	when	"01101010",	--(X"8")	106
          "10011001"	when	"01101011",	--(X"99")	107
          "10001011"	when	"01101100",	--(X"8b")	108
          "00011101"	when	"01101101",	--(X"1d")	109
          "11110010"	when	"01101110",	--(X"f2")	110
          "10110100"	when	"01101111",	--(X"b4")	111
          "11101001"	when	"01110000",	--(X"e9")	112
          "11000111"	when	"01110001",	--(X"c7")	113
          "10011111"	when	"01110010",	--(X"9f")	114
          "01001010"	when	"01110011",	--(X"4a")	115
          "00110001"	when	"01110100",	--(X"31")	116
          "00100101"	when	"01110101",	--(X"25")	117
          "11111110"	when	"01110110",	--(X"fe")	118
          "01111100"	when	"01110111",	--(X"7c")	119
          "11010011"	when	"01111000",	--(X"d3")	120
          "10100010"	when	"01111001",	--(X"a2")	121
          "10111101"	when	"01111010",	--(X"bd")	122
          "01010110"	when	"01111011",	--(X"56")	123
          "00010100"	when	"01111100",	--(X"14")	124
          "10001000"	when	"01111101",	--(X"88")	125
          "01100000"	when	"01111110",	--(X"60")	126
          "00001011"	when	"01111111",	--(X"0b")	127
          "11001101"	when	"10000000",	--(X"cd")	128
          "11100010"	when	"10000001",	--(X"e2")	129
          "00110100"	when	"10000010",	--(X"34")	130
          "01010000"	when	"10000011",	--(X"50")	131
          "10011110"	when	"10000100",	--(X"9e")	132
          "11011100"	when	"10000101",	--(X"dc")	133
          "00010001"	when	"10000110",	--(X"11")	134
          "00000101"	when	"10000111",	--(X"5")	135
          "00101011"	when	"10001000",	--(X"2b")	136
          "10110111"	when	"10001001",	--(X"b7")	137
          "10101001"	when	"10001010",	--(X"a9")	138
          "01001000"	when	"10001011",	--(X"48")	139
          "11111111"	when	"10001100",	--(X"ff")	140
          "01100110"	when	"10001101",	--(X"66")	141
          "10001010"	when	"10001110",	--(X"8a")	142
          "01110011"	when	"10001111",	--(X"73")	143
          "00000011"	when	"10010000",	--(X"3")	144
          "01110101"	when	"10010001",	--(X"75")	145
          "10000110"	when	"10010010",	--(X"86")	146
          "11110001"	when	"10010011",	--(X"f1")	147
          "01101010"	when	"10010100",	--(X"6a")	148
          "10100111"	when	"10010101",	--(X"a7")	149
          "01000000"	when	"10010110",	--(X"40")	150
          "11000010"	when	"10010111",	--(X"c2")	151
          "10111001"	when	"10011000",	--(X"b9")	152
          "00101100"	when	"10011001",	--(X"2c")	153
          "11011011"	when	"10011010",	--(X"db")	154
          "00011111"	when	"10011011",	--(X"1f")	155
          "01011000"	when	"10011100",	--(X"58")	156
          "10010100"	when	"10011101",	--(X"94")	157
          "00111110"	when	"10011110",	--(X"3e")	158
          "11101101"	when	"10011111",	--(X"ed")	159
          "11111100"	when	"10100000",	--(X"fc")	160
          "00011011"	when	"10100001",	--(X"1b")	161
          "10100000"	when	"10100010",	--(X"a0")	162
          "00000100"	when	"10100011",	--(X"4")	163
          "10111000"	when	"10100100",	--(X"b8")	164
          "10001101"	when	"10100101",	--(X"8d")	165
          "11100110"	when	"10100110",	--(X"e6")	166
          "01011001"	when	"10100111",	--(X"59")	167
          "01100010"	when	"10101000",	--(X"62")	168
          "10010011"	when	"10101001",	--(X"93")	169
          "00110101"	when	"10101010",	--(X"35")	170
          "01111110"	when	"10101011",	--(X"7e")	171
          "11001010"	when	"10101100",	--(X"ca")	172
          "00100001"	when	"10101101",	--(X"21")	173
          "11011111"	when	"10101110",	--(X"df")	174
          "01000111"	when	"10101111",	--(X"47")	175
          "00010101"	when	"10110000",	--(X"15")	176
          "11110011"	when	"10110001",	--(X"f3")	177
          "10111010"	when	"10110010",	--(X"ba")	178
          "01111111"	when	"10110011",	--(X"7f")	179
          "10100110"	when	"10110100",	--(X"a6")	180
          "01101001"	when	"10110101",	--(X"69")	181
          "11001000"	when	"10110110",	--(X"c8")	182
          "01001101"	when	"10110111",	--(X"4d")	183
          "10000111"	when	"10111000",	--(X"87")	184
          "00111011"	when	"10111001",	--(X"3b")	185
          "10011100"	when	"10111010",	--(X"9c")	186
          "00000001"	when	"10111011",	--(X"1")	187
          "11100000"	when	"10111100",	--(X"e0")	188
          "11011110"	when	"10111101",	--(X"de")	189
          "00100100"	when	"10111110",	--(X"24")	190
          "01010010"	when	"10111111",	--(X"52")	191
          "01111011"	when	"11000000",	--(X"7b")	192
          "00001100"	when	"11000001",	--(X"0c")	193
          "01101000"	when	"11000010",	--(X"68")	194
          "00011110"	when	"11000011",	--(X"1e")	195
          "10000000"	when	"11000100",	--(X"80")	196
          "10110010"	when	"11000101",	--(X"b2")	197
          "01011010"	when	"11000110",	--(X"5a")	198
          "11100111"	when	"11000111",	--(X"e7")	199
          "10101101"	when	"11001000",	--(X"ad")	200
          "11010101"	when	"11001001",	--(X"d5")	201
          "00100011"	when	"11001010",	--(X"23")	202
          "11110100"	when	"11001011",	--(X"f4")	203
          "01000110"	when	"11001100",	--(X"46")	204
          "00111111"	when	"11001101",	--(X"3f")	205
          "10010001"	when	"11001110",	--(X"91")	206
          "11001001"	when	"11001111",	--(X"c9")	207
          "01101110"	when	"11010000",	--(X"6e")	208
          "10000100"	when	"11010001",	--(X"84")	209
          "01110010"	when	"11010010",	--(X"72")	210
          "10111011"	when	"11010011",	--(X"bb")	211
          "00001101"	when	"11010100",	--(X"0d")	212
          "00011000"	when	"11010101",	--(X"18")	213
          "11011001"	when	"11010110",	--(X"d9")	214
          "10010110"	when	"11010111",	--(X"96")	215
          "11110000"	when	"11011000",	--(X"f0")	216
          "01011111"	when	"11011001",	--(X"5f")	217
          "01000001"	when	"11011010",	--(X"41")	218
          "10101100"	when	"11011011",	--(X"ac")	219
          "00100111"	when	"11011100",	--(X"27")	220
          "11000101"	when	"11011101",	--(X"c5")	221
          "11100011"	when	"11011110",	--(X"e3")	222
          "00111010"	when	"11011111",	--(X"3a")	223
          "10000001"	when	"11100000",	--(X"81")	224
          "01101111"	when	"11100001",	--(X"6f")	225
          "00000111"	when	"11100010",	--(X"7")	226
          "10100011"	when	"11100011",	--(X"a3")	227
          "01111001"	when	"11100100",	--(X"79")	228
          "11110110"	when	"11100101",	--(X"f6")	229
          "00101101"	when	"11100110",	--(X"2d")	230
          "00111000"	when	"11100111",	--(X"38")	231
          "00011010"	when	"11101000",	--(X"1a")	232
          "01000100"	when	"11101001",	--(X"44")	233
          "01011110"	when	"11101010",	--(X"5e")	234
          "10110101"	when	"11101011",	--(X"b5")	235
          "11010010"	when	"11101100",	--(X"d2")	236
          "11101100"	when	"11101101",	--(X"ec")	237
          "11001011"	when	"11101110",	--(X"cb")	238
          "10010000"	when	"11101111",	--(X"90")	239
          "10011010"	when	"11110000",	--(X"9a")	240
          "00110110"	when	"11110001",	--(X"36")	241
          "11100101"	when	"11110010",	--(X"e5")	242
          "00101001"	when	"11110011",	--(X"29")	243
          "11000011"	when	"11110100",	--(X"c3")	244
          "01001111"	when	"11110101",	--(X"4f")	245
          "10101011"	when	"11110110",	--(X"ab")	246
          "01100100"	when	"11110111",	--(X"64")	247
          "01010001"	when	"11111000",	--(X"51")	248
          "11111000"	when	"11111001",	--(X"f8")	249
          "00010000"	when	"11111010",	--(X"10")	250
          "11010111"	when	"11111011",	--(X"d7")	251
          "10111100"	when	"11111100",	--(X"bc")	252
          "00000010"	when	"11111101",	--(X"2")	253
          "01111101"	when	"11111110",	--(X"7d")	254
          "10001110"	when	"11111111",	--(X"8e")	255           
                                                         
         "XXXXXXXX" WHEN OTHERS;

end Behavioral;
